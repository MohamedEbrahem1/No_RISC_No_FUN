`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/06/2023 11:40:32 AM
// Design Name: 
// Module Name: jump_ctrl
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module jump_generator(
input [1:0] jump,
input [9:0] PC,
input [31:0] result,
output reg [31:0] jump_result
    );
        
endmodule
